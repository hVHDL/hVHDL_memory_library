
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package dual_port_ram_pkg is

    constant read_pipeline_delay : natural := 2;
    type ram_array is array (natural range <>) of std_logic_vector;

    type ram_in_record is record
        address           : unsigned;
        read_is_requested : std_logic;
        data              : std_logic_vector;
        write_requested   : std_logic;
    end record;

    type ram_out_record is record
        data          : std_logic_vector;
        data_is_ready : std_logic;
    end record;

    type ram_in_array is array (natural range <>) of ram_in_record;
    type ram_out_array is array (natural range <>) of ram_out_record;

    type dpram_ref_record is record
        ram_in       : ram_in_record;
        ram_out      : ram_out_record;
        address_high : natural;
        data         : std_logic_vector;
        address      : std_logic_vector;
    end record;

    function create_ref_subtypes(datawidth : natural; addresswidth : natural) return dpram_ref_record;

    procedure init_ram (
        signal self_in : out ram_in_record);

    procedure init_ram (
        signal self_in : inout ram_in_array);

    procedure request_data_from_ram (
        signal self_in : out ram_in_record;
        address : in natural);

    function ram_read_is_ready ( self_read_out : ram_out_record)
        return boolean;

    function get_ram_data ( self_read_out : ram_out_record)
        return std_logic_vector;

    function get_uint_ram_data ( self_read_out : ram_out_record)
        return integer;
------------------------------------------------------------------------
------------------------------------------------------------------------
    procedure write_data_to_ram (
        signal self_in : out ram_in_record;
        address : in natural;
        data    : in std_logic_vector);

    function write_requested_to_address(ram_in : ram_in_record; address : natural) 
        return boolean;

end package dual_port_ram_pkg;

package body dual_port_ram_pkg is

------------------------------------------------------------------------
    function create_ref_subtypes(datawidth : natural; addresswidth : natural) return dpram_ref_record is
        constant retval : dpram_ref_record :=
        (
            ram_in => (
                address            => (0 to addresswidth-1  => '0')
                ,read_is_requested => '0'
                ,data              => (datawidth-1 downto 0 => '0')
                ,write_requested   => '0')

            ,ram_out =>(
                data           => (datawidth-1 downto 0 => '0')
                ,data_is_ready => '0')
            
            ,address_high => 2**addresswidth - 1
            ,data    => (datawidth-1 downto 0    => '0')
            ,address => (addresswidth-1 downto 0 => '0')
        );
    begin
        return retval;
    end create_ref_subtypes;
------------------------------------------------------------------------
    procedure init_ram
    (
        signal self_in : out ram_in_record
    ) is
    begin
        self_in.read_is_requested <= '0';
        self_in.write_requested   <= '0';
    end init_ram;

    procedure init_ram
    (
        signal self_in : inout ram_in_array
    ) is
    begin
        for i in self_in'range loop
            self_in(i).read_is_requested <= '0';
            self_in(i).write_requested <= '0';
        end loop;
    end init_ram;

------------------------------
    procedure request_data_from_ram
    (
        signal self_in : out ram_in_record;
        address : in natural
    ) is
    begin

        self_in.address <= to_unsigned(address, self_in.address'length);
        self_in.read_is_requested <= '1';

    end request_data_from_ram;
------------------------------
    function ram_read_is_ready
    (
        self_read_out : ram_out_record
    )
    return boolean
    is
    begin
        return self_read_out.data_is_ready = '1';
        
    end ram_read_is_ready;
------------------------------
    function get_ram_data
    (
        self_read_out : ram_out_record
    )
    return std_logic_vector 
    is
    begin
        return self_read_out.data;
    end get_ram_data;
------------------------------------------------------------------------
    function get_uint_ram_data
    (
        self_read_out : ram_out_record
    )
    return integer
    is
    begin
        return to_integer(unsigned(self_read_out.data));
    end get_uint_ram_data;
------------------------------------------------------------------------
------------------------------------------------------------------------
    procedure write_data_to_ram
    (
        signal self_in : out ram_in_record;
        address : in natural;
        data : in std_logic_vector
    ) is
    begin
        self_in.address <= to_unsigned(address, self_in.address'length);
        self_in.data    <= data;
        self_in.write_requested <= '1';
    end write_data_to_ram;
------------------------------------------------------------------------
    function write_requested_to_address(ram_in : ram_in_record; address : natural) return boolean is
    begin
        return ram_in.write_requested = '1' and ram_in.address = address;
    end write_requested_to_address;
------------------------------------------------------------------------
end package body dual_port_ram_pkg;
------------------------------------------------------------------------
------------------------------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

    use work.dual_port_ram_pkg.all;

entity dual_port_ram is
    generic(
       g_dpram_subtype : dpram_ref_record
       ; g_ram_init_values : work.dual_port_ram_pkg.ram_array
           (0 to g_dpram_subtype.address_high
           )(
           g_dpram_subtype.data'range) := (others => (others => '0')));

    port (
        clock     : in std_logic;
        ram_a_in  : in work.dual_port_ram_pkg.ram_in_record;
        ram_a_out : out work.dual_port_ram_pkg.ram_out_record;
        --------------------
        ram_b_in  : in work.dual_port_ram_pkg.ram_in_record;
        ram_b_out : out work.dual_port_ram_pkg.ram_out_record
    );
end entity dual_port_ram;
