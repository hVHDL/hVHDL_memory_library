library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;

package fpga_dual_port_ram_pkg is

end package fpga_dual_port_ram_pkg;

package body fpga_dual_port_ram_pkg is

end package body fpga_dual_port_ram_pkg;
